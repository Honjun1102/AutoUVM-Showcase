`ifndef AUTOUVM_CLK_RST_IF_SV
`define AUTOUVM_CLK_RST_IF_SV

interface autouvm_clk_rst_if;
    logic clk;
    logic rst;
endinterface

`endif
