// AutoUVM自动生成 - AXI4 Sequencer

class cpu_axi4_sequencer extends uvm_sequencer #(axi4_transaction);
  `uvm_component_utils(cpu_axi4_sequencer)
  
  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction
  
endclass
